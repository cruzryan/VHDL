library IEEE;

use IEEE.std_logic_1164.ALL;

ENTITY EAPriory is

	PORT(
		I: IN STD_LOGIC_VECTOR(8 downto 0);
        DISPLAY: OUT STD_LOGIC_VECTOR(6 downto 0)
		);

end EAPriory;

ARCHITECTURE main of EAPriory IS
BEGIN
	PROCESS
	BEGIN

	CASE I IS
		WHEN "000000000" => DISPLAY <= "0000001";
		WHEN "100000000" => DISPLAY <= "1001111";
		WHEN "110000000" => DISPLAY <= "0010010";
		WHEN "111000000" => DISPLAY <= "0000110";
		WHEN "111100000" => DISPLAY <= "1001101";
		WHEN "111110000" => DISPLAY <= "0100100";
		WHEN "111111000" => DISPLAY <= "1100000";
		WHEN "111111100" => DISPLAY <= "0001111";
		WHEN "111111110" => DISPLAY <= "0000000";
		WHEN OTHERS => DISPLAY <= "0001100";
	END CASE;

	wait for 10 ns;
	END PROCESS;
end ARCHITECTURE;